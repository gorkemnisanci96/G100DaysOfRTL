// Clock Gating Levels
//1- Gating the clock at the source level. 
//2-Gating the clock in the module level 
//3-Gating the clock in the flop level 
